`timescale 1ns / 1ps
//////////////////////////////////////////////////////////////////////////////////
// Company: 
// Engineer: 
// 
// Create Date:    19:18:39 11/11/2015 
// Design Name: 
// Module Name:    Seg7_Dev 
// Project Name: 
// Target Devices: 
// Tool versions: 
// Description: 
//
// Dependencies: 
//
// Revision: 
// Revision 0.01 - File Created
// Additional Comments: 
//
//////////////////////////////////////////////////////////////////////////////////
module Seg7_Dev(
    input [2:0]Scan,
    input [31:0]Hexs,
    input flash_clk,
    input [7:0]point,
    input [7:0]LES,
    output [7:0]SEGMENT,
    output [3:0]AN
    );


endmodule
