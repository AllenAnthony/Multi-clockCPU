`timescale 1ns / 1ps
//////////////////////////////////////////////////////////////////////////////////
// Company: 
// Engineer: 
// 
// Create Date:    19:09:12 11/11/2015 
// Design Name: 
// Module Name:    InputT32 
// Project Name: 
// Target Devices: 
// Tool versions: 
// Description: 
//
// Dependencies: 
//
// Revision: 
// Revision 0.01 - File Created
// Additional Comments: 
//
//////////////////////////////////////////////////////////////////////////////////
module InputT32(
    input [2:0]push_out,
    input [4:0]disp_ctr,
    output [31:0]Ai,
    output [31:0]Bi,
    output [1:0]state,
    output [3:0]blink
    );


endmodule
